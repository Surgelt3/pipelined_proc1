module extend(input [31:7] instr,
                input [1:0] immsrc,
                output reg [31:0] immext);
    
    always @(*) begin

        case (immsrc)
            // i type instrucitions
            2'b00: immext = {{20{instr[31]}}, instr[31:20]};

            // s type
            2'b01: immext = {{20{instr[31]}}, instr[31:25], instr[11:7]};
            //b type
            2'b10: immext = {{20{instr[31]}}, instr[31:20]};
            // jtype
            2'b11: immext = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};

            default: immext = 32'bx;
    
        endcase

    end



endmodule